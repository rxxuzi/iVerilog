module COMP_EQ(a,b,a_eq_b);
input a,b;
output a_eq_b;

assign a_eq_b= (a==b);

endmodule

