// コメントのテスト
/* コメントのテスト */
module gand(a,b,c);     
input a,b;
output c;
assign c=a&b;     // コメントのテスト
endmodule
